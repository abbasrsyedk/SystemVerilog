interface intf(input logic clk,reset);
  
  //declaring the signals
  logic       en;
  logic [3:0] count_out;
  
endinterface