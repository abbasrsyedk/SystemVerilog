interface mux_intf();
	logic x;
	logic y;
    logic z;
    logic m;
    logic [1:0]select;
	logic mux_out;
endinterface
